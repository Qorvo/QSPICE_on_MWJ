* QSPICE_on_MWJ\Article4\Sim1\VRM_PSRR_OnOff.qsch
Rload VOUT 0 100
Vac N05 N01 AC 1
Vref REF 0 DC 0.5
Vin N01 0 DC 10
M_PMOS VOUT N02 VIN VIN PFET PMOS
Cout N03 N04 22µ
Rfb VOUT FB 90K
Rg FB 0 10K
Copen N07 0 {Copen}
L1 N08 N07 {Lopen}
EA N06 0 FB REF 3K
Vsine VIN N05 SIN 0 1m 10Meg
R2 VOUT N03 10m
L2 N04 0 1n
Rbw N06 N08 1Meg
Cbw N08 0 22p
Ebuf N02 0 N07 0 1
.model PFET PMOS Kp=100 eta=10m VT0 = -1
.param Lopen={if(x, 1f, 1K)}
.param Copen={if(x, 1f, 1K)}
.step param x list 0 1
.ac dec 20 1 100Meg
.plot AC 1/V(VOUT)
.lib PMOS.txt
.end
