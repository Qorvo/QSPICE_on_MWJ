* C:\Users\mn080015\OneDrive - Qorvo\Documents\QSPICE\QSPICE_on_MWJ_SIJ\Article3\Sim1\VRM_PSRR_LineReg_sch.qsch
Rload VOUT 0 100
Vripple VIN N04 AC 1
Vref N08 0 DC 0.5
Vin N04 0 DC 10
�1 N01 N02 N10 N07 N03 � � � � � � � � � � � RRopAmp Avol=20 GBW=47Meg Slew=100Meg Rload=10 Phi=90
V15 N01 0 15
Vm15 N02 0 -15
M_PMOS VOUT N09 VIN VIN PFET PMOS
Cout N11 N06 47�
Resr VOUT N11 1m
Lesl N06 0 0.2n
Rfb VOUT N03 90K
Rg N03 0 10K
Elinereg N05 N08 VIN N08 0.2m
Rnr N05 N07 1Meg
Cnr N07 0 10n
Lopen N10 N09 {L_open}
Copen N09 0 {C_open}
.model PFET PMOS Kp=1000 eta=10m
.ac dec 10 1 10Meg
.plot AC 1/V(VOUT)
.param L_open={if(x, 1f, 1K)}
.param C_open={if(x, 1f, 1K)}
.step param x list 0 1
.lib PMOS.txt
.end
