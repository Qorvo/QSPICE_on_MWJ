* C:\Users\mn080015\OneDrive - Qorvo\Documents\QSPICE\QSPICE_on_MWJ_SIJ\Article2\Sim2\VRM_PSRR.qsch
Rload VOUT 0 100
Vripple VIN N04 AC 1
Vref N09 0 DC 0.5
Vin N04 0 DC 10
�1 N01 N02 N07 N09 N03 � � � � � � � � � � � RRopAmp Avol=20 GBW=47Meg Slew=100Meg Rload=10 Phi=90
V15 N01 0 15
Vm15 N02 0 -15
M_PMOS VOUT N06 VIN VIN PFET PMOS
Cout N08 N05 47�
Resr VOUT N08 1m
Lesl N05 0 0.2n
Rfb VOUT N03 90K
Rg N03 0 10K
Lopen N07 N06 {L_open}
Copen N06 0 {C_open}
.model PFET PMOS Kp=1000 eta=10m
.ac dec 10 1 10Meg
.plot AC 1/V(VOUT)
.param L_open={if(x, 1f, 1K)}
.param C_open={if(x, 1f, 1K)}
.step param x list 0 1
.lib PMOS.txt
.end
