* C:\Users\mn080015\OneDrive - Qorvo\Documents\QSPICE\QSPICE_on_MWJ_SIJ\Article2\Sim1\VRM_GainBW.qsch
Rload VOUT 0 100
Vac N07 N06 AC 1
Vref N06 0 DC 0.5
Vin VIN 0 DC 10
�1 N01 N02 N05 N07 N03 � � � � � � � � � � � RRopAmp Avol=20 GBW=47Meg Slew=100Meg Rload=10 Phi=90
V15 N01 0 15
Vm15 N02 0 -15
M_PMOS VOUT N05 VIN VIN PFET PMOS
Cout VOUT 0 47�
Rfb VOUT N04 90K
Rg N04 0 10K
Lopen N03 N04 {L_open}
Copen N03 0 {C_open}
.model PFET PMOS Kp=1000 eta=10m
.ac dec 10 1 10Meg
.plot AC V(VOUT)
.param L_open={if(x, 1f, 1K)}
.param C_open={if(x, 1f, 1K)}
.step param x list 0 1
.lib PMOS.txt
.end
