* QSPICE_on_MWJ\Article2\Sim1\VRM_GainBW.qsch
Rload VOUT 0 {Rload}
Vac N07 N06 AC 1
Vref N06 0 DC 0.5
Vin VIN 0 DC 10
M_PMOS VOUT N02 VIN VIN PFET PMOS
Cout N03 0 22�
Rfb VOUT N01 90K
Rg N01 0 10K
Copen FB 0 {Copen}
L1 FB N01 {Lopen}
EA N04 0 FB REF 3K
Vsine REF N07 SIN 0 1m 100K
R2 VOUT N03 10m
Rbw N04 N05 1Meg
Cbw N05 0 22p
Ebuf N02 0 N05 0 1
.model PFET PMOS Kp=100 eta=10m VT0 = -1
.param Lopen={if(x, 1f, 1K)}
.param Copen={if(x, 1f, 1K)}
.step param x list 0 1
.param Rload 100
.ac dec 20 1 100Meg
.plot AC V(VOUT)
*.param Rload 1
*.tran 100�
*.plot tran V(VOUT)
.lib PMOS.txt
.end
